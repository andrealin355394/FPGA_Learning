`timescale 1ns/1ns
module tb ();








initial #1000 $stop;  // modelsim simulator stop condition
                      // don't delete
endmodule
